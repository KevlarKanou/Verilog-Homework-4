module tb (

);

endmodule